----------------------------------------------------------------------------------
-- Create Date                       : 09/19/2016 10:30:22 AM
-- Module Name                       : fft_engine - Behavioral
-- company                           : Airbus Group India Pvt.Ltd
-- Engineer                          : Vishal Goyal, Sourabh Tapas
-- Development Platform              : Vivado 2016.1
-- Testing and Verification Platform : Vivado 2016.1
-- Target Devices                    : KC705 Evaluation Board for the Kintex-7 FPGA
------------------------------------------------------------------------------------

library ieee;
library unisim;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use unisim.vcomponents.all;
use ieee.std_logic_signed.all;

entity fft_engine is
port ( clk_primary_p        : in  std_logic;                                                                -- Primary system clock input
       clk_primary_n        : in  std_logic;                                                                -- - LVDS.
        
       clk_10               : out std_logic;                                                                -- 10 Mhz Clock.
       cpi_trigger          : in  std_logic;                                                                -- Coherent pulse interval trigger.
       rst                  : in  std_logic;                                                                -- Active high reset - synchronous to clock.
       rd_en                : in  std_logic;                                                                -- Read enable. Used by external master(previous module) to signal that it is able to provide meaningful data.
       num_of_samples       : in  std_logic_vector( 7 downto 0);                                            -- Length/number of samples(payload size) defined by user [ configurable value can be anything between decimal(0 to 61) ]
       dpc_fft_Im           : in  std_logic_vector(15 downto 0);                                            -- Inphase/real part of Input channel. Carries the unprocessed sample data: XN_RE.
       dpc_fft_Qm           : in  std_logic_vector(15 downto 0);                                            -- Quadraturephase/imaginary part of Input channel. Carries the unprocessed sample data: XN_IM.
       wr_en                : out std_logic;                                                                -- Write Enable. Generated by the fft IP core to signal that it is able to provide processed sample data.
       s_axis_data_tready   : out std_logic;                                                                -- TREADY for the Data Input channel. Generated by the fft core to signal that it is ready to accept data.
       fft_cfar_Im          : out std_logic_vector(15 downto 0);                                            -- Inphase/real part of fft engine's output channel.Carries the processed sample data: XK_RE.
       fft_cfar_Qm          : out std_logic_vector(15 downto 0);                                            -- Quadraturephase/imaginary part of fft engine's output channel.Carries the processed sample data: XK_IM.
       doppler_cell         : out std_logic_vector( 5 downto 0);                                            -- FFT core output sample index on the scale of 0 to 63 in natural order. 
       cnt63_pin            : out std_logic_vector( 7 downto 0));                                           -- Decimal 64 counter.
end fft_engine;

architecture Behavioral of fft_engine is

-- component declaration of clock wizard IP - generated by the Clocking Wizard

component CLK_wiz
port( clk_primary_p  : in std_logic;
      clk_primary_n  : in std_logic;                                                                       
      clk_10         : out std_logic);                                                                     
end component;

-- ccmponent declaration of metastability hardener for the incoming reset

component meta_harden is
Port ( clk_dst    : in  std_logic;
       rst_dst    : in  std_logic;
       signal_src : in  std_logic;
       signal_dst : out std_logic);
end component meta_harden;

-- 64 points Fast Fourier Transform IP component Declaration

component fft_IP 
port ( 
  -- General signals
       aclk                        : in  std_logic;                                                        -- Rising-edge clock
       aclken                      : in  std_logic;                                                        -- Active-High clock enable (optional)
       aresetn                     : in  std_logic;                                                        -- Active-Low synchronous clear (optional, always take priority over aclken) A minimum aresetn active pulse of two cycles is required.

  -- Config slave channel signals        
       s_axis_config_tdata         : in  std_logic_vector(7 downto 0);                                     -- TDATA  for the Configuration channel. Carries the configuration information: CP_LEN, FWD/INV,NFFT and SCALE_SCH.
       s_axis_config_tvalid        : in  std_logic;                                                        -- TVALID for the Configuration channel. Asserted by the external master to signal that it is able to provide data.
       s_axis_config_tready        : out std_logic;                                                        -- TREADY for the Configuration channel. Asserted by the core to signal that it is ready to accept data.
  
  -- Data slave channel signals  
       s_axis_data_tdata           : in  std_logic_vector(31 downto 0);                                    -- TDATA  for the Data Input channel. Carries the unprocessed sample data: XN_RE and XN_IM.
       s_axis_data_tvalid          : in  std_logic;                                                        -- TVALID for the Data Input channel. Used by the external master to signal that it is able to provide data.
       s_axis_data_tready          : out std_logic;                                                        -- TREADY for the Data Input channel. Used by the core to signal that it is ready to accept data.
       s_axis_data_tlast           : in  std_logic;                                                        -- TLAST  for the Data Input channel. Asserted by the external master on the last sample of the frame. This is not used by the core except to generate the events event_tlast_unexpected and event_tlast_missing events.

  -- Data master channel signals
       m_axis_data_tdata           : out std_logic_vector(31 downto 0);                                    -- TDATA  for the Data Output channel. Carries the processed sample data XK_RE and XK_IM
       m_axis_data_tuser           : out std_logic_vector(7 downto 0);                                     -- TUSER  for the Data Output channel. Carries additional per-sample information, such as XK_INDEX, OVFLO and BLK_EXP.
       m_axis_data_tvalid          : out std_logic;                                                        -- TVALID for the Data Output channel. Asserted by the core to signal that it is able to provide sample data.
       m_axis_data_tready          : in  std_logic;                                                        -- TREADY for the Data Output channel. Asserted by the external slave to signal that it is ready to accept data. Only present in "Non-Realtime" mode.
       m_axis_data_tlast           : out std_logic;                                                        -- TLAST  for the Data Output channel. Asserted by the core on the last sample of the frame.

  -- Event signals
       event_frame_started         : out std_logic;                                                        -- Asserted when the core starts to process a new frame.
       event_tlast_unexpected      : out std_logic;                                                        -- Asserted when the core sees s_axis_data_tlast High on a data sample that is not the last one in a frame.
       event_tlast_missing         : out std_logic;                                                        -- Asserted when s_axis_data_tlast is Low on the last data sample of a frame.
       event_status_channel_halt   : out std_logic;                                                        -- Asserted when the core tries to write data to the Status channel and it is unable to do so. Only present in "Non-Realtime" mode.
       event_data_in_channel_halt  : out std_logic;                                                        -- Asserted when the core requests data from the Data Input channel and none is available.
       event_data_out_channel_halt : out std_logic);                                                       -- Asserted when the core tries to write data to the Data Output channel and it is unable to do so. Only present in "Non-Realtime" mode.
end component;

-- signal declaration
    -- Memory generator signals

        signal rangecell                   : integer range 0 to 1670:= 0;                                  -- Rangecell count (incerments after each frame of 64 samples)
        signal cnt63                       : std_logic_vector(7 downto 0);                                 -- Decimal 64 counter.
        signal clk_10_s, not_rst,rst_s     : std_logic;                                                    -- 10 Mhz clock signal for intermididate operations, inverted reset signal and metahardened reset signal.


    -- fft portmap signals
    
        signal s_axis_data_tlast_s         : std_logic;                                                    -- TLAST signal for the Data Input channel
        signal s_axis_data_tready_s        : std_logic;                                                    -- TREADY for the Data Input channel. Used by the fft core to signal that it is ready to accept data.
        signal s_axis_config_tdata_s       : std_logic_vector(7 downto 0):= "00000001";                    -- TDATA  for the Configuration channel. Carries the configuration information: CP_LEN, FWD/INV,NFFT and SCALE_SCH.
        signal dpc_fft_Im_s                : std_logic_vector(15 downto 0);                                -- Inphase/real part of Input channel.  Carries the unprocessed sample data: XN_RE.
        signal dpc_fft_Qm_s                : std_logic_vector(15 downto 0);                                -- Quadraturephase/imaginary part of Input channel.Carries the unprocessed sample data: XN_IM. 
        signal doppler_cell_s              : std_logic_vector(7 downto 0);
        
begin

-- signal connections

not_rst            <= not rst;                                                                             -- Generating active low reset signal for fft IP 
clk_10             <= clk_10_s;                                                                            -- Connect 10 MHz clock signal to 10 MHz clock port pin
cnt63_pin          <= cnt63;                                                                               -- Connect decimal 64 count to count 64 pin 
doppler_cell       <= doppler_cell_s(5 downto 0);                                                          -- Connect doppler cell signal with doppler cell port
s_axis_data_tready <= s_axis_data_tready_s;                                                                -- Connect s_axis_data_tready_s signal to s_axis_data_tready port

-- Component Instantiations

FFT_IP_inst: fft_IP 
port map ( aclk                            => clk_10_s,
           aclken                          => '1',
           aresetn                         => not_rst,
           ---------------------------------------------------------
           s_axis_config_tdata             => s_axis_config_tdata_s,
           s_axis_config_tvalid            => '1',
           s_axis_config_tready            => open,
           ----------------------------------------------------------
           s_axis_data_tdata(15 downto 0)  => dpc_fft_Im_s,
           s_axis_data_tdata(31 downto 16) => dpc_fft_Qm_s,
           s_axis_data_tvalid              => rd_en,
           s_axis_data_tready              => s_axis_data_tready_s,
           s_axis_data_tlast               => s_axis_data_tlast_s,
           ---------------------------------------------------------
           m_axis_data_tdata(15 downto 0)  => fft_cfar_Im,
           m_axis_data_tdata(31 downto 16) => fft_cfar_Qm,
           m_axis_data_tuser               => doppler_cell_s,
           m_axis_data_tvalid              => wr_en,
           m_axis_data_tready              => '1',                                                          -- This pin can be taken out as port in entity if needed as control signal to make connection with next module CFAR.
           m_axis_data_tlast               => open,
           ---------------------------------------------------------
           event_frame_started             => open,
           event_tlast_unexpected          => open,
           event_tlast_missing             => open,
           event_status_channel_halt       => open,
           event_data_in_channel_halt      => open,
           event_data_out_channel_halt     => open);

Clock_wizard_inst: CLK_wiz
port map ( clk_primary_p => clk_primary_p,
           clk_primary_n => clk_primary_n,
           clk_10        => clk_10_s);
           
meta_hard_rst: meta_harden
port map ( rst_dst    => '0',
           clk_dst    => clk_10_s,
           signal_src => rst, 
           signal_dst => rst_s);

-----------------------------------------------------------------------------------------------------------

-- Zero_padding

    dpc_fft_Im_s <=  dpc_fft_Im when cnt63 >= 2 and cnt63 <= (num_of_samples + 2) else (others => '0');    -- padding enough number of zero samples to make payload sample length to 64 samples for Im
    dpc_fft_Qm_s <=  dpc_fft_Qm when cnt63 >= 2 and cnt63 <= (num_of_samples + 2) else (others => '0');    -- padding enough number of zero samples to make payload sample length to 64 samples for Qm
                                                                                                           -- +2 is done because to take care of Latency from BROM 
-- tlast signal generation

    s_axis_data_tlast_s <= '1' when cnt63 = "00111111" else '0';                                           -- makimg tlast signal high for 1 clock cycle on last sample of 64 point size fft 

-- Decimal 64 counter 

sample_cnt_64:process(clk_10_s)
begin 
    if rising_edge(clk_10_s) then                                                                          -- synchronous event test
        if(rst_s = '1') then                                                                               -- Reset synchronous to clock
            cnt63 <= (others => '0');                                                                      -- reset the counter
            rangecell <= 0;                                                                                -- reset the rangecell
        else                                                                                               -- non-reset behavior
            if rd_en = '1' and s_axis_data_tready_s = '1' then                                             -- Checking, whether fft_engine ready to accept data and external device providing valid data?
                if rangecell < 1667 then                                                                   -- Yes, then check is rangecell count is less than 1667?
                    if (cnt63 < 63) then                                                                   -- Yes, then check is count63 is less than 63?
                       cnt63 <= cnt63 + '1';                                                               -- Yes, then increment count63 by 1
                    else                                                                                   -- No, then
                        cnt63    <= (others => '0');                                                       -- reinitialise the count to zero
                        rangecell <= rangecell + 1;                                                        -- increment the rangecell
                    end if;                                                                                -- end of cnt63 condition
                else                                                                                       -- rangecell is not less than 1667 then
                    rangecell <= 0;                                                                        -- reinitialise the rangecell to zero
                    cnt63 <= cnt63 + '1';                                                                  -- increment count63 by 1
                end if;                                                                                    -- end of rangecell condition
            else                                                                                           -- fft_engine is not ready to accept the data or external device is not providing valid data yet then
                cnt63    <= (others => '0');                                                               -- reset the counter
            end if;                                                                                        -- end of ready signal checking condition
        end if;                                                                                            -- end of reset/normal operation
    end if;                                                                                                -- end of synchronous events
end process;
end Behavioral;