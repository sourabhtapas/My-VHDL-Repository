----------------------------------------------------------------------------------
-- Create Date                       : 04/08/2016 12:27:16 PM
-- Module Name                       : Digital Pulse Compression Block (DPC)
-- company                           : Airbus Group India Pvt.Ltd
-- Engineer                          : Vishal Goyal, Sourabh Tapas
-- Development Platform              : Vivado 2016.1
-- Testing and Verification Platform : Vivado 2016.1
----------------------------------------------------------------------------------

library ieee;
library unisim;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;
use unisim.vcomponents.all;
use work.all;
use work.mydatatype_pkg.all;                                   -- To load P2 code and P4 code coefficients

entity DPC_module is
Port ( dpc_clk_in_p    : in  std_logic;                        -- primary system clock input
       dpc_clk_in_n    : in  std_logic;                        -- - LVDS
       clk5            : out std_logic;                        -- 5 MHz clock
       clk30           : out std_logic;                        -- 30 MHz clock
       locked          : out std_logic;                        -- locked of clock wizard
       rst             : in  std_logic;                        -- active high reset - synchronous to clock
       I_main          : in  std_logic_vector (15 downto 0);   -- Input  correspoding to Inphase part of Main channel
       Q_main          : in  std_logic_vector (15 downto 0);   -- Input  correspoding to Quadraturephase part of Main channel
       I_aux           : in  std_logic_vector (15 downto 0);   -- Input  correspoding to Inphase part of Auxilary channel
       Q_aux           : in  std_logic_vector (15 downto 0);   -- Input  correspoding to Quadraturephase part of Auxilary channel
       dpcOut_Imain16  : out std_logic_vector (15 downto 0);   -- Output correspoding to Inphase part of Main channel
       dpcOut_Qmain16  : out std_logic_vector (15 downto 0);   -- Output correspoding to Quadraturephase part of Main channel
       dpcOut_Iaux16   : out std_logic_vector (15 downto 0);   -- Output correspoding to Inphase part of Auxilary channel
       dpcOut_Qaux16   : out std_logic_vector (15 downto 0));  -- Output correspoding to Quadraturephase part of Auxilary channel
end DPC_module; 


architecture Behavioral of DPC_module is

-- creating memory of size: width = 16 and depth = 196 

Type sr196X16 is array (0 to 195) of std_logic_vector (15 downto 0);
signal a, b, f, g : sr196X16;                                       -- memory arrays for tapped delay line structure 


-- Internal signals

signal s_coef                                                      : aslv98X17;                          -- multiplexed signal to feed data of six channels one by one on rotation basis to Mul_Acc component
signal s_pair                                                      : aslv98X18;                          -- multiplexed signal to feed data of six channels one by one on rotation basis to Mul_Acc component
signal clk5_s, clk30_s, locked_s                                   : std_logic;                          -- 5 MHz clock,30 MHz clock, locked of clock wizard and active high reset respectively
signal a_pair,aplusb_pair,bsuba_pair,f_pair,fplusg_pair,gsubf_pair : aslv98X18;                          -- memory array signals to store folded input data
signal CS                                                          : std_logic_vector (2  downto 0);     -- channel select (CS) 3 bit counter signal
signal p, s, w, t, r, v                                            : std_logic_vector (35 downto 0);     -- Demultiplexed signals from Mul_Acc output one by one on rotation basis
signal dpcOut_Imain, dpcOut_Qmain, dpcOut_Iaux, dpcOut_Qaux        : std_logic_vector (35 downto 0);     -- memory signal to store FIR structure's final output at every rising edge of 5 MHz clock
signal A_out0_s, A_out1_s, A_out2_s, A_out3_s, A_out4_s, A_out5_s  : std_logic_vector (35 downto 0);     -- signals to connect with Mul_Acc Component


-- ccmponent declaration of clock wizard IP - generated by the Clocking Wizard

component CLK_Wiz
port( clk_in1_p  : in  std_logic;
      clk_in1_n  : in  std_logic;
      clk_out_30 : out std_logic;
      clk_out_5  : out std_logic;
      locked     : out std_logic);
end component;


-- ccmponent declaration of metastability hardener for the incoming reset

--component meta_harden is
--Port ( clk_dst    : in  std_logic;
--       rst_dst    : in  std_logic;
--       signal_src : in  std_logic;
--       signal_dst : out std_logic);
--end component meta_harden;


-- component declaration of Mul_Acc

component Mul_Acc
Port ( CLK          : in  std_logic;
       coef         : in  aslv98X17;
       pair         : in  aslv98X18;
       reset        : in  std_logic;
       A_out0       : out std_logic_vector (35 downto 0);
       A_out1       : out std_logic_vector (35 downto 0);
       A_out2       : out std_logic_vector (35 downto 0);
       A_out3       : out std_logic_vector (35 downto 0);
       A_out4       : out std_logic_vector (35 downto 0);
       A_out5       : out std_logic_vector (35 downto 0));
end component;


begin

clk5 <= clk5_s;                                            -- Connect 5 MHz clock signal to 5 MHz clock port pin
clk30 <= clk30_s;                                          -- Connect 30 MHz clock signal to 30 MHz clock port pin
locked <= locked_s;                                        -- Connect locked signal of clock wizard to locked port pin


-- Instantiate clk_core 

CLK_IP: CLK_Wiz
port map ( clk_in1_p  => dpc_clk_in_p,
           clk_in1_n  => dpc_clk_in_n,
           clk_out_30 => clk30_s,
           clk_out_5  => clk5_s,
           locked     => locked_s);
           
-- Instantiate a metastability hardener for the incoming reset

--meta_hard_rst: meta_harden
--port map ( rst_dst    => '0',
--           clk_dst    => clk5_s,
--           signal_src => rst, 
--           signal_dst => rst_s);


-- Tapped delay line structure/shift register structure  for Imain, Qmain, Iauxilary and Qauxilary channels.

Delay_line: process(clk5_s)
    begin
        if(rising_edge(clk5_s)) then                                               -- synchronous event test
            if (rst = '1') then                                                    -- active high reset - synchronous to clock
                a <= (others =>(others=>'0')); b <= (others =>(others=>'0'));      -- clear all the memory data when reset condition is true (high)
                f <= (others =>(others=>'0')); g <= (others =>(others=>'0'));
            else                                                                   -- non-reset behavior
                a(0) <= I_main;  a(1 to 195) <=  a(0 to 194);                      -- New data enters on 0th location and  
                b(0) <= Q_main;  b(1 to 195) <=  b(0 to 194);                      -- - previous data is shifted to the next location on every rising edge of 5 MHz clock
                f(0) <= I_aux;   f(1 to 195) <=  f(0 to 194);                      -- - for each memory array (i.e for a,b,f,g)
                g(0) <= Q_aux;   g(1 to 195) <=  g(0 to 194);
            end if;                                                                -- end of reset/normal operation
        end if;                                                                    -- end of synchronous events
end process Delay_line;


-- As the codes are a lot symmetric we half the number of multiplier by folding the FIR structure so that one multiplier gets addition of two inputs
-- ( refer last but one paragraph on 1st page of "Digital Pulse Compression Block.docx" for clarification )

a_pair_set: for i in 0 to 97 generate
begin
    a_pair(i) <= (((a(i)(15)&a(i)(15)&a(i)(15 downto 0)) + ((a(195 - i)(15)&a(195 - i)(15)&a(195 - i)(15 downto 0)))));        -- for P2 code
                
end generate;

aplusb_pair_set: for i in 0 to 97 generate
begin
    aplusb_pair(i) <= (((a(i)(15)&a(i)(15)&a(i)(15 downto 0)) + ((a(195 - i)(15)&a(195 - i)(15)&a(195 - i)(15 downto 0)))) + ((b(i)(15)&b(i)(15)&b(i)(15 downto 0)) + ((b(195 - i)(15)&b(195 - i)(15)&b(195 - i)(15 downto 0)))));              -- for P2 code
                     
end generate;

bsuba_pair_set: for i in 0 to 97 generate
begin
    bsuba_pair(i) <= (((b(i)(15)&b(i)(15)&b(i)(15 downto 0)) + ((b(195 - i)(15)&b(195 - i)(15) & b(195 - i)(15 downto 0)))) - ((a(i)(15)&a(i)(15)&a(i)(15 downto 0)) + ((a(195 - i)(15)&a(195 - i)(15)&a(195 - i)(15 downto 0)))));             -- for P2 code
                     
end generate;

f_pair_set: for i in 0 to 97 generate
begin
    f_pair(i) <= (((f(i)(15)&f(i)(15)&f(i)(15 downto 0)) + ((f(195 - i)(15)&f(195 - i)(15)&f(195 - i)(15 downto 0))))) ;        -- for P2 code
                 
end generate;

fplusg_pair_set: for i in 0 to 97 generate
begin
    fplusg_pair(i) <= (((f(i)(15)&f(i)(15)&f(i)(15 downto 0)) + ((f(195 - i)(15)&f(195 - i)(15)&f(195 - i)(15 downto 0)))) + ((g(i)(15)&g(i)(15)&g(i)(15 downto 0)) + ((g(195 - i)(15)&g(195 - i)(15)&g(195 - i)(15 downto 0)))));        -- for P2 code
                      
end generate;

gsubf_pair_set: for i in 0 to 97 generate
begin
    gsubf_pair(i) <= (((g(i)(15)&g(i)(15)&g(i)(15 downto 0)) + ((g(195 - i)(15)&g(195 - i)(15)&g(195 - i)(15 downto 0)))) - ((f(i)(15)&f(i)(15)&f(i)(15 downto 0)) + ((f(195 - i)(15)&f(195 - i)(15)&f(195 - i)(15 downto 0)))));              -- for P2 code
                     
end generate;


--free running counter of decimal 6 to detect rising edge of 30 MHz clock.

ch_select: process(clk30_s)
begin
    if rising_edge(clk30_s) then          -- synchronous event test
        if(rst = '1') then                -- active high reset - synchronous to clock
            CS  <= "000";                 -- reset the counter
        else                              -- non-reset behavior
            if (CS = "101") then          -- Is count equal to "101"?
                CS <= "000";              -- Yes, then reset the count to all zero
            else                          -- No, 
                CS  <= CS + 1;            -- then Increment the count by 1
            end if;                       -- end of counter condition
        end if;                           -- end of reset/normal operation
    end if;                               -- end of synchronous events
end process ch_select;


-- multiplexing and Demultiplexing of signal to to Mul_Acc component for six channels one by one on rotation basis

Channel_wheel: process(CS, a_pair, f_pair, aplusb_pair, fplusg_pair, bsuba_pair, gsubf_pair, A_out0_s, A_out1_s, A_out2_s, A_out3_s, A_out4_s, A_out5_s)
begin
case CS is
when "000" =>

            s_coef  <=  P2_coefCplusD;                           -- for P4 code
            s_pair  <=  a_pair;
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
when "001" =>

            s_coef  <=  P2_coefCplusD;                           -- for P2 code
            s_pair  <=  f_pair;
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
when "010" =>

            s_coef  <=  P2_coefD;                                -- for P2 code
            s_pair  <=  aplusb_pair;
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
when "011" =>
 
            s_coef  <=  P2_coefD;                                -- for P2 code
            s_pair  <=  fplusg_pair;
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
when "100" =>

                s_coef  <=  P2_coefC;                                -- for P2 code

            s_pair  <=  bsuba_pair;
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
when "101" =>

            s_coef  <=  P2_coefC;                           -- for P2 code
            s_pair  <=  gsubf_pair;
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
when others =>
            s_coef  <=  p2_coefCplusD;                           -- any value, it doesn't matter 
            s_pair  <=  a_pair;                                  -- any value, it doesn't matter 
            p       <=  A_out0_s;
            s       <=  A_out1_s;
            w       <=  A_out2_s;
            t       <=  A_out3_s;
            r       <=  A_out4_s;
            v       <=  A_out5_s;
end case;
end process;


-- Instantiation of Mul_Acc component ( Multiplier and Accumulator )

MAC: Mul_Acc
port map ( CLK    => clk30_s,
           coef   => s_coef,
           pair   => s_pair,
           reset  => rst,               
           A_out0 => A_out0_s,
           A_out1 => A_out1_s,
           A_out2 => A_out2_s,
           A_out3 => A_out3_s,
           A_out4 => A_out4_s, 
           A_out5 => A_out5_s);


-- Final Output of DPC Module

Output: process(clk5_s)
begin
   if(rising_edge(clk5_s)) then                                                        -- synchronous event test
       if rst = '1' then                                                               -- active high reset - synchronous to clock
                dpcOut_Imain <= (others => '0');   dpcOut_Qmain <= (others => '0');
                dpcOut_Iaux  <= (others => '0');   dpcOut_Qaux  <= (others => '0');    -- clear all the outputs when reset condition is true (high)
            else                                                                       -- non-reset behavior
                dpcOut_Imain <= ((p) - (w));   dpcOut_Qmain <= ((p) + (r));            -- refer 1st page of "Digital Pulse Compression Block.docx"  (p - w) is equivalent to (K1- K2) and (p + r) is equivalent to (K1 + K3) for Main channel output
                dpcOut_Iaux  <= ((s) - (t));   dpcOut_Qaux  <= ((s) + (v));            -- refer 1st page of "Digital Pulse Compression Block.docx"  (s - t) is equivalent to (K1- K2) and (s + v) is equivalent to (K1 + K3) for Auxilary Channel output
       end if;                                                                         -- end of reset/normal operation
   end if;                                                                             -- end of synchronous events
end process Output;
                dpcOut_Imain16 <= dpcOut_Imain(35 downto 20);                          -- resizing Actual 36 bit output to 16 bit   
                dpcOut_Qmain16 <= dpcOut_Qmain(35 downto 20);                          -- resizing Actual 36 bit output to 16 bit
                dpcOut_Iaux16  <= dpcOut_Iaux (35 downto 20);                          -- resizing Actual 36 bit output to 16 bit 
                dpcOut_Qaux16  <= dpcOut_Qaux (35 downto 20);                          -- resizing Actual 36 bit output to 16 bit 
end Behavioral;