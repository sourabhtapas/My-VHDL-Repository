----------------------------------------------------------------------------------
-- Create Date                       : 09/19/2016 10:30:22 AM
-- Module Name                       : hw_env_fft - Behavioral
-- company                           : Airbus Group India Pvt.Ltd
-- Engineer                          : Vishal Goyal, Sourabh Tapas
-- Development Platform              : Vivado 2016.1
-- Testing and Verification Platform : Vivado 2016.1
-- Target Devices                    : KC705 Evaluation Board for the Kintex-7 FPGA
----------------------------------------------------------------------------------

library ieee;
library unisim;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use unisim.vcomponents.all;
use ieee.std_logic_signed.all;

entity hw_env_fft is
port ( clk_primary_p           : in  std_logic;                                                             -- primary system clock input
       clk_primary_n           : in  std_logic;                                                             -- - LVDS
       hw_rst                  : in  std_logic;                                                             -- active high reset - synchronous to clock
       hw_fft_cfar_Im          : out std_logic_vector(15 downto 0);                                         -- Inphase/real part of fft engine's output channel.Carries the processed sample data: XK_RE.
       hw_fft_cfar_Qm          : out std_logic_vector(15 downto 0));                                        -- Quadraturephase/imaginary part of fft engine's output channel.Carries the processed sample data: XK_IM.
end hw_env_fft;

architecture Behavioral of hw_env_fft is

component fft_engine
port ( clk_primary_p        : in  std_logic;                                                                -- Primary system clock input
       clk_primary_n        : in  std_logic;                                                                -- - LVDS.
        
       clk_10               : out std_logic;                                                                -- 10 Mhz Clock.
       cpi_trigger          : in  std_logic;                                                                -- Coherent pulse interval trigger.
       rst                  : in  std_logic;                                                                -- Active high reset - synchronous to clock.
       rd_en                : in  std_logic;                                                                -- Read enable. Used by external master(previous module) to signal that it is able to provide meaningful data.
       num_of_samples       : in  std_logic_vector( 7 downto 0);                                            -- Length/number of samples(payload size) defined by user [ configurable value can be anything between decimal(0 to 61) ]
       dpc_fft_Im           : in  std_logic_vector(15 downto 0);                                            -- Inphase/real part of Input channel. Carries the unprocessed sample data: XN_RE.
       dpc_fft_Qm           : in  std_logic_vector(15 downto 0);                                            -- Quadraturephase/imaginary part of Input channel. Carries the unprocessed sample data: XN_IM.
       wr_en                : out std_logic;                                                                -- Write Enable. Generated by the fft IP core to signal that it is able to provide processed sample data.
       s_axis_data_tready   : out std_logic;                                                                -- TREADY for the Data Input channel. Generated by the fft core to signal that it is ready to accept data.
       fft_cfar_Im          : out std_logic_vector(15 downto 0);                                            -- Inphase/real part of fft engine's output channel.Carries the processed sample data: XK_RE.
       fft_cfar_Qm          : out std_logic_vector(15 downto 0);                                            -- Quadraturephase/imaginary part of fft engine's output channel.Carries the processed sample data: XK_IM.
       doppler_cell         : out std_logic_vector( 5 downto 0);                                            -- FFT core output sample index on the scale of 0 to 63 in natural order. 
       cnt63_pin            : out std_logic_vector( 7 downto 0));                                           -- Decimal 64 counter.
end component;

component BROM_Im
port ( clka  : in std_logic;
       ena   : in std_logic;
       addra : in std_logic_vector(16 downto 0);
       douta : out std_logic_vector(15 downto 0));
end component;

component BROM_Qm
port ( clka  : in std_logic;
       ena   : in std_logic;
       addra : in std_logic_vector(16 downto 0);
       douta : out std_logic_vector(15 downto 0));
end component;

component BROM_Im_1
port ( clka  : in std_logic;
       ena   : in std_logic;
       addra : in std_logic_vector(16 downto 0);
       douta : out std_logic_vector(15 downto 0));
end component;

component BROM_Qm_1
port ( clka  : in std_logic;
       ena   : in std_logic;
       addra : in std_logic_vector(16 downto 0);
       douta : out std_logic_vector(15 downto 0));
end component;        

-- signal declaration

        signal rd_addr_slv                                            : std_logic_vector(16 downto 0);     -- Read address counter for Input data memory location address in standard logic vector data type
        signal rd_addr                                                : integer range 0 to 106690 := 0;    -- Read address counter for Input data memory location address
        signal ptr                                                    : integer range 0 to 106690 := 0;    -- Pointer register as counter for the generation of CPI_trigger signal
        signal s_axis_data_tready_s                                   : std_logic;                         -- TREADY for the Data Input channel. Used by the fft core to signal that it is ready to accept data
        signal clk_10_s                                               : std_logic;                         -- 10 Mhz clock signal 
        signal rd_en_s                                                : std_logic := '0';                  -- Read enable signal as a tready signal for the Data Input channel
        signal cpi_trigger_s                                          : std_logic:= '0';                   -- Coherent pulse interval trigger signal
        signal toggle                                                 : std_logic := '0';                  -- Select input of multiplexer to switch between test vector sets/two data bursts
        signal dpc_data_Im, dpc_data_Qm, dpc_data_Im_1, dpc_data_Qm_1 : std_logic_vector(15 downto 0);     -- Multiplexed input data channels of respective test vector set
        signal dpc_in_Im, dpc_in_Qm                                   : std_logic_vector(15 downto 0);     -- Multiplexed output data channel of multiplexer
        signal cnt63                                                  : std_logic_vector(7 downto 0);      -- Decimal 64 counter 
        signal num_of_samples_s                                       : std_logic_vector(7 downto 0);      -- Configurable user defined value of length/number of samples( payload size) coming from previous DPC module

begin

fft_engine_inst: fft_engine  
port map ( clk_primary_p                   => clk_primary_p,
           clk_primary_n                   => clk_primary_n,
           
           s_axis_data_tready              => s_axis_data_tready_s,
           cpi_trigger                     => cpi_trigger_s,
           clk_10                          => clk_10_s,
           rst                             => hw_rst,
           rd_en                           => rd_en_s,
           dpc_fft_Im                      => dpc_in_Im,
           dpc_fft_Qm                      => dpc_in_Qm,
           wr_en                           => open,
           fft_cfar_Im                     => hw_fft_cfar_Im,  
           fft_cfar_Qm                     => hw_fft_cfar_Qm,
           num_of_samples                  => num_of_samples_s,
           doppler_cell                    => open,
           cnt63_pin                       => cnt63);           

BROM_Imain_inst: BROM_Im
port map ( clka  => clk_10_s,
           ena   => '1',
           addra => rd_addr_slv,
           douta => dpc_data_Im);

BROM_Imain_1_inst: BROM_Im_1
port map ( clka  => clk_10_s,
           ena   => '1',
           addra => rd_addr_slv,
           douta => dpc_data_Im_1);          
          
BROM_Qmain_inst: BROM_Qm
port map ( clka  => clk_10_s,
           ena   => '1',
           addra => rd_addr_slv,
           douta => dpc_data_Qm);

BROM_Qmain_1_inst: BROM_Qm_1
port map ( clka  => clk_10_s,
           ena   => '1',
           addra => rd_addr_slv,
           douta => dpc_data_Qm_1);

-- test vector Selection

    dpc_in_Im <= dpc_data_Im when toggle = '0' else dpc_data_Im_1;                                         -- Multiplexer to switch between test vector sets for Im
    dpc_in_Qm <= dpc_data_Qm when toggle = '0' else dpc_data_Qm_1;                                         -- Multiplexer to switch between test vector sets for Qm

-- Data address generations and synchronised tunning


Read_address: process(clk_10_s)
begin
   if rising_edge(clk_10_s) then                                                                           -- Synchronous event test
       if(hw_rst = '1') then                                                                               -- Reset synchronous to clock
           rd_addr <= 0;                                                                                   -- Reset the rd_addr counter
       else                                                                                                -- Non-reset behavior
           if rd_en_s = '1' and s_axis_data_tready_s = '1' then                                            -- Checking, whether fft_engine ready to accept data and whether external device providing valid data?
               if (rd_addr < (("0000011010000011")*(num_of_samples_s + '1'))) then                         -- Yes, then check is read address less than for e.g.80016 (for 48 samples)? [ 1667 X 48 = 80016 is the total number of samples in first test vector set when toggle = 0][ 1667 X 50 = 83350 is the total number of samples in second test vector when toggle = 1]. "0000011010000011" is binary equivalent of 1667. This conversion is required because data type should be same for multiply operation. 
                   if (cnt63 <= num_of_samples_s) then                                                     -- Yes, then check is cnt63 less than num_of_samples(i.e. user defined payload size)?
                       rd_addr <= rd_addr + 1;                                                             -- Yes, then increment the reading address
                   else                                                                                    -- No, then
                           rd_addr <= rd_addr;                                                             -- Hold the read address value
                   end if;                                                                                 -- End of cnt63 check condition
               else                                                                                        -- Read address is not less than 80016 then
                   rd_addr <= 0;                                                                           -- Re-initialise the address to zero 
               end if;                                                                                     -- End of read address counter condition
           end if;                                                                                         -- End of ready signal checking condition
       end if;                                                                                             -- End of reset/normal operation
   end if;                                                                                                 -- End of synchronous events
end process read_address;

rd_addr_slv <= std_logic_vector(to_unsigned(rd_addr,rd_addr_slv'length));                                  -- Converting decimal rd_addr to standard logic vector data type

-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- Generation of control signals
-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
CPI_trigger_generation: process(clk_10_s)
begin
    if rising_edge(clk_10_s) then                                                                           -- Synchronous event test
       if(hw_rst = '1') then                                                                                -- reset synchronous to clock
             ptr <= 106670;                                                                                 -- Reset the pointer value to 106670 (  Any value can be taken ) [ chosen just to witness qucker generation of cpi_trigger initially ]
        else                                                                                                -- Non-reset behavior       
            if (ptr < 106687) then                                                                          -- Is pointer less than 106687? [ 1667 X 64 = 106688 is the total number of samples after doing the zero padding to 48 input damples ]  
                ptr <= ptr + 1;                                                                             -- Yes, then increment the pointer   
            else                                                                                            -- Pointer is not less than 106687                  
                ptr  <= 0;                                                                                  -- Then re-initialise the pointer to zero
            end if;                                                                                         -- End of pointer counter condition
        end if;                                                                                             -- End of reset/normal operation
    end if;                                                                                                 -- End of synchronous events
end process;


    cpi_trigger_s    <= '1'        when ptr = 106687 else '0';                                              -- Generation of CPI_trigger pulse after every burst[ i.e. after 1667 X 64 = 106688 samples].

    num_of_samples_s <= "00101111" when toggle = '0' else "00110001";                                       -- Assigning user defined value say 47(i.e.48 sample payload size) first and say 49( i.e.50 sample payload size) on next burst to show configurable feature of FFT_engine module
    
rd_pro: process(cpi_trigger_s)
begin 
    if (cpi_trigger_s = '1') then
      rd_en_s <= '1';                                                                                       -- Generation of read enable as soon as first cpi_trigger arrives to indicate that valid data is available from previous module (i.e.DPC)
    end if;
end process;

    -- switching of test vector at cpi_trigger event
        
        switch_tvec_at_cpi: process(clk_10_s)
        begin 
            if rising_edge(clk_10_s) then                                                                                   -- Synchronous event test
                if (cpi_trigger_s = '1') then -- OR -- if (rising_edge(cpi_trigger_s) then (will also work on ILA)          -- Is cpi_trigger high?
                    toggle <= not toggle;                                                                                   -- Yes, then invert the toggle signal and hold till next cpi_trigger pulse arrives
                end if;                                                                                                     -- End of cpi_trigger check condition
            end if;                                                                                                         -- End of synchronous events
        end process;

-- Known issue:
-- Below line/ lines of code is/are equivalent of above switch_tvec_at_cpi process and gives exactly same clean waveforms in Behavioral simulation but for no real reason on Kintex FPGA kit (as shown by waveforms in ILA)the
-- toggle signal errorneously inverting before last but one rangecell of burst causing missing of last rangecell data and duplication of next burst's first rangecell data in it's place.

--    toggle      <= not toggle when rising_edge(cpi_trigger_s);
    
                  -- OR --

-- switch_tvec_at_cpi: process(cpi_trigger_s)
--            begin 
--                if rising_edge(cpi_trigger_s) then                                                           -- Is cpi_trigger high?
--                    toggle <= not toggle;                                                                    -- Yes, then invert the toggle signal and hold till next cpi_trigger pulse arrives
--                end if;                                                                                      -- End of cpi_trigger check condition
--            end process;

end Behavioral;